///////////////////////////////////////////////////////
parameter NOP = 32'b0000000_00000_00000_00000_0000000000; //NOP
parameter ADD = 32'b0000010_00001_00010_00011_0000000000; // Add	r1,r2,r3 //4110C00
parameter SUB = 32'b0000101_00100_00001_00011_0000000000; // Sub	r4,r1,r3 //A408C00
parameter SLT = 32'b1100101_00001_00010_00011_0000000000; // slt	if R2 < R3 then R1 = 1
parameter AND = 32'b0001000_00001_00010_00011_0000000000; // AND: R1 <- R2 AND R3
parameter OR =  32'b0001010_00001_00010_00011_0000000000; // OR:  R1 <- R2 OR R3
parameter XOR = 32'b0001100_00001_00010_00011_0000000000; // XOR: R1 <- R2 XOR R3
parameter ST =  32'b0000001_00000_00100_00001_0000000000; // ST:  M[R4] <- R1
parameter LD =  32'b0100001_00100_00001_00000_0000000000; // LD:  R1 <- M[R4]
parameter ADI = 32'b0100010_00001_00010_000000000000001; // ADI: R1 <- R2 + 1 
parameter SBI = 32'b0100101_00001_00010_000000000000001; // SBI: R1 <- R2 - 1
parameter NOT = 32'b0101110_00001_00010_000000000000000; // NOT: R1 <- ~R2 
parameter ANI = 32'b0101000_00001_00010_000000000000001; // ANI: R1 <- R2 AND 000...1
parameter ORI = 32'b0101010_00001_00010_000000000000000; // ORI: R1 <- R2 OR  000...0
parameter XRI = 32'b0101100_00001_00010_000000000000000; // XRI: R1 <- R2 XOR 000...0
parameter AIU = 32'b1100010_00001_00010_000000000000001; // AIU: R1 <- R2 + 1
parameter SIU = 32'b1000101_00001_00010_000000000000001; // SIU: R1 <- R2 - 1
parameter MOV = 32'b1000000_00011_00001_000000000000000; // MOV: R1 <- R3
parameter LSL = 32'b0110000_00001_00010_000000000000001; // LSL: R1 <- R2 << 1
parameter LSR = 32'b0110001_00001_00010_000000000000001; // LSR: R1 <- R2 >> 1
parameter ASL = 32'b0110010_00001_00010_000000000000001; // ASL: R1 <- R2 <<< 1
parameter ASR = 32'b0110011_00001_00010_000000000000001; // ASR: R1 <- R2 >>> 1
parameter ROL = 32'b0110100_00001_00010_000000000000001; // ROL: R1 <- {R2[30:0],R2[31]}
parameter ROR = 32'b0110101_00001_00010_000000000000001; // ROR: R1 <- {R2[0],R2[31:1]}
parameter JMR = 32'b1100001_00000_00010_000000000000000; // JMR: PC <- R0
parameter BZ =  32'b0100000_00000_00010_000000000000001; // BZ:  if R0=0 PC <- (PC+1)+1
parameter BNZ = 32'b1100000_00000_00010_000000000000001; // BNZ: if R0!=0 PC <- (PC+1)+1
parameter JMP = 32'b1000100_00000_00010_000000000000001; // JMP: PC <- (PC+1)+1
parameter JML = 32'b0000111_00001_00010_000000000000000; // JML: PC <- (PC+1)+1, R1 <- PC+1
///////////////////////////////////////////////////////





